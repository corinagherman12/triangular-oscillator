** Profile: "SCHEMATIC1-bias"  [ C:\Users\corin\OneDrive\Desktop\P1\SIMULARE\simulare-pspicefiles\schematic1\bias.sim ] 

** Creating circuit file "bias.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "C:/Users/corin/OneDrive/Desktop/P1/biblioteci spice/bc846b.lib" 
.LIB "C:/Users/corin/OneDrive/Desktop/P1/biblioteci spice/bc856b.lib" 
.LIB "C:/Users/corin/OneDrive/Desktop/P1/biblioteci spice/bzx84c2v7.lib" 
.LIB "C:/Users/corin/OneDrive/Desktop/P1/biblioteci spice/diode.lib" 
* From [PSPICE NETLIST] section of C:\Users\corin\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 10ms 100u 1u SKIPBP 
.TEMP 0,30,70
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
